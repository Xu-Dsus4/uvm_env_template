`include "ut/xsc_test/env/seq_lib/xsc_sequence0.svh"